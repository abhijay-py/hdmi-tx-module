
module hdmi_tx_top (
    input logic clk, n_rst,
    output logic hdmi_clk_p, hdmi_clk_n, hdmi_hpd, hdmi_scl, hdmi_sda, hdmi_cec
    output logic [2:0] hdmi_p, hdmi_n
)


endmodule